module  vv(
i,
o,
o1
);

input i;
output reg o=i;
output reg o1;

endmodule 
