
 module  i1  
  
 (
      );
 input     a  ;
 
 output     b  ;
 
 output     c  ;
 
 assign        b  =  ( 1 +  ( 2 + 1 )  * 3 * 4 )  +  ( 1 +  ( 2 + 1 )  + 3 * 4 )  + 3 * 4 - 1 +  ( 2 + 1 )  + 1 +  ( 2 + 1 )  + 3 * 4 ;
 
 assign        c  = 7 - 5 + 1 ;
 
 
 endmodule
 