`line 1 src/define.v 1
`line 3 src/define.v 1

`line 5 src/define.v 1
`line 6 src/define.v 1
`line 9 src/define.v 1
`line 12 src/define.v 1
module i1();

input a;
output b;
output c;
assign b = (1+(2+1)*3* 4)+(1+(2+1)+3* 4) +3* 4-1+(2+1) + 1+(2+1) +3* 4 ;
assign c = 7-  
  5 + 
	
12 +
21 +1;

endmodule


