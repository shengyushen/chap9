
 module  ssy  
  
 (
      );
 parameter    p1  = 1121 ;
 
 integer  i1  = 1345 ;
 
 integer  i2  = 4'b11_00 ;
 
 integer  i3  = 4'd1122 ;
 
 integer  i4  = 4'h11_22 ;
 
 integer  i5  = 4'o11_22 ;
 
 
 endmodule
 