module empty();
endmodule



