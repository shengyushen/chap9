module ssy();
parameter p1 = 11_21;
integer i1= 13_45;
integer i2 = 4'b11_00;
integer i3 = 4'D11_22;
integer i4 = 4'h11_22;
integer i5 = 4'O11_22;
endmodule
