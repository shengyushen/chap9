module i1();

endmodule
//sdf
