
module xx();
output gg;
assign gg=    1 +   2 ;
endmodule

