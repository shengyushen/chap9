module test;
	parameter x = "String with escaped backslash at end \\";
	initial
		$display("PASSED");
endmodule
