module t(
	input a ,
	output b
);

assign b = 1;


endmodule


`line 1 ./src/test_step2_define.v 1 






module i(input a,b,c,output o2,o3);
assign o2 = a+b;
assign o3 = a+b+ c;

endmodule

`line 14 src/test_step2_reverse_define.v 2 

