
       module    i1    
       (        )  ;     
 endmodule
   